
// a class is a dynamic object and a module is a static object 
// so when we say static we mean that when we performe a simulation the module object will be there right from the start of our simulation tell the end even if we do not use it
// Whereas when we consider a class, we may require to use an object from a class and when we no longer need it we could just delete it during a simulation.
class first;                         
                                      
  reg [2:0] data; 
  reg [1:0] data2;
  
  
endclass
 
 
module tb;
  
  first f;
  
  initial begin
    f = new();// here we use new in order to create an object which means that we are allocating a memory for our object
              //if we don't do it f object will be just a NULL pointer
    f.data = 3'b111;// here is how we can access the atributs of our object
    f.data2 = 2'b01;
    
    f = null;// here we deallocate the memory of our object means f will be pointing to null again
    
    #1;
    $display("Value of data : %0d and data2 : %0d",f.data, f.data2);
  end
  
  
  
endmodule

 // if we use a module instead of class  in verilog
/*====================================*/
module top( input a, b, output y);
  reg temp;
  assign y = a & b; // this a continous assignment
  
endmodule

//we use the module here

module top2(input c, d, output e);
  
  top dut(c, d, e);// this is how we create an instance of our module
  dut.temp; // here is how to access a variable of our object
  
endmodule

/*===================================*/



// in general functions are just like in c language 
module test();
  
  // we could also initialize the arguments in function declaration
  /* we could use add() as folow
  function bit[7:0] add();
  
    return a + b;
  
  endfunction
  -> but in this case a and b should be visible to the function 
  
  ===============================================
  or we could also use the following declaration
  
  function void add(input bit[6:0] a, b);
  
    $display("a = %0d and b = %0d ", a, b);
    
  
  endfunction
  
  -> we refere to this declaration in case we want to display variables or somthing
  ================================================
  we can not controling time using a function 
  because time controling is not allowed inside a function
  for that we use task  instead
  */
  function bit[7:0] add(input bit[6:0] a, b);
  
    return a + b;
  
  endfunction
  
  bit [6:0] ain = 3, bin = 6;

  bit[9:0] res = 0;

  initial begin
	// we could do this 
    res = add(4, 3);
    // we could also do this 
    res = add(ain, bin);
    // and this
    res = add(); /* but in this case we have declare "a" and "b" before declaring the 							function so that they will be visible to the add function*/
    $display("result is -> %0d", res);

  end
    
endmodule
